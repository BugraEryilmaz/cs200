module dpiempty();
    export "DPI-C" function tmp;
    function tmp();
    endfunction
endmodule